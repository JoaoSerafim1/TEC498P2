module tablememory7by5 (
cell0_0S, cell1_0S, cell2_0S, cell3_0S, cell4_0S, cell5_0S, cell6_0S,
cell0_1S, cell1_1S, cell2_1S, cell3_1S, cell4_1S, cell5_1S, cell6_1S,
cell0_2S, cell1_2S, cell2_2S, cell3_2S, cell4_2S, cell5_2S, cell6_2S,
cell0_3S, cell1_3S, cell2_3S, cell3_3S, cell4_3S, cell5_3S, cell6_3S,
cell0_4S, cell1_4S, cell2_4S, cell3_4S, cell4_4S, cell5_4S, cell6_4S,

cell0_0R, cell1_0R, cell2_0R, cell3_0R, cell4_0R, cell5_0R, cell6_0R,
cell0_1R, cell1_1R, cell2_1R, cell3_1R, cell4_1R, cell5_1R, cell6_1R,
cell0_2R, cell1_2R, cell2_2R, cell3_2R, cell4_2R, cell5_2R, cell6_2R,
cell0_3R, cell1_3R, cell2_3R, cell3_3R, cell4_3R, cell5_3R, cell6_3R,
cell0_4R, cell1_4R, cell2_4R, cell3_4R, cell4_4R, cell5_4R, cell6_4R,

cell0_0Q, cell1_0Q, cell2_0Q, cell3_0Q, cell4_0Q, cell5_0Q, cell6_0Q,
cell0_1Q, cell1_1Q, cell2_1Q, cell3_1Q, cell4_1Q, cell5_1Q, cell6_1Q,
cell0_2Q, cell1_2Q, cell2_2Q, cell3_2Q, cell4_2Q, cell5_2Q, cell6_2Q,
cell0_3Q, cell1_3Q, cell2_3Q, cell3_3Q, cell4_3Q, cell5_3Q, cell6_3Q,
cell0_4Q, cell1_4Q, cell2_4Q, cell3_4Q, cell4_4Q, cell5_4Q, cell6_4Q
);

	input
	cell0_0S, cell1_0S, cell2_0S, cell3_0S, cell4_0S, cell5_0S, cell6_0S,
	cell0_1S, cell1_1S, cell2_1S, cell3_1S, cell4_1S, cell5_1S, cell6_1S,
	cell0_2S, cell1_2S, cell2_2S, cell3_2S, cell4_2S, cell5_2S, cell6_2S,
	cell0_3S, cell1_3S, cell2_3S, cell3_3S, cell4_3S, cell5_3S, cell6_3S,
	cell0_4S, cell1_4S, cell2_4S, cell3_4S, cell4_4S, cell5_4S, cell6_4S,

	cell0_0R, cell1_0R, cell2_0R, cell3_0R, cell4_0R, cell5_0R, cell6_0R,
	cell0_1R, cell1_1R, cell2_1R, cell3_1R, cell4_1R, cell5_1R, cell6_1R,
	cell0_2R, cell1_2R, cell2_2R, cell3_2R, cell4_2R, cell5_2R, cell6_2R,
	cell0_3R, cell1_3R, cell2_3R, cell3_3R, cell4_3R, cell5_3R, cell6_3R,
	cell0_4R, cell1_4R, cell2_4R, cell3_4R, cell4_4R, cell5_4R, cell6_4R;
	
	output
	cell0_0Q, cell1_0Q, cell2_0Q, cell3_0Q, cell4_0Q, cell5_0Q, cell6_0Q,
	cell0_1Q, cell1_1Q, cell2_1Q, cell3_1Q, cell4_1Q, cell5_1Q, cell6_1Q,
	cell0_2Q, cell1_2Q, cell2_2Q, cell3_2Q, cell4_2Q, cell5_2Q, cell6_2Q,
	cell0_3Q, cell1_3Q, cell2_3Q, cell3_3Q, cell4_3Q, cell5_3Q, cell6_3Q,
	cell0_4Q, cell1_4Q, cell2_4Q, cell3_4Q, cell4_4Q, cell5_4Q, cell6_4Q;

srlt_gate cell0_0 (
		.q (cell0_0Q),
		.s (cell0_0S),
		.r (cell0_0R)
);

srlt_gate cell1_0 (
		.q (cell1_0Q),
		.s (cell1_0S),
		.r (cell1_0R)
);

srlt_gate cell2_0 (
		.q (cell2_0Q),
		.s (cell2_0S),
		.r (cell2_0R)
);

srlt_gate cell3_0 (
		.q (cell3_0Q),
		.s (cell3_0S),
		.r (cell3_0R)
);

srlt_gate cell4_0 (
		.q (cell4_0Q),
		.s (cell4_0S),
		.r (cell4_0R)
);

srlt_gate cell5_0 (
		.q (cell5_0Q),
		.s (cell5_0S),
		.r (cell5_0R)
);

srlt_gate cell6_0 (
		.q (cell6_0Q),
		.s (cell6_0S),
		.r (cell6_0R)
);

srlt_gate cell0_1 (
		.q (cell0_1Q),
		.s (cell0_1S),
		.r (cell0_1R)
);

srlt_gate cell1_1 (
		.q (cell1_1Q),
		.s (cell1_1S),
		.r (cell1_1R)
);

srlt_gate cell2_1 (
		.q (cell2_1Q),
		.s (cell2_1S),
		.r (cell2_1R)
);

srlt_gate cell3_1 (
		.q (cell3_1Q),
		.s (cell3_1S),
		.r (cell3_1R)
);

srlt_gate cell4_1 (
		.q (cell4_1Q),
		.s (cell4_1S),
		.r (cell4_1R)
);

srlt_gate cell5_1 (
		.q (cell5_1Q),
		.s (cell5_1S),
		.r (cell5_1R)
);

srlt_gate cell6_1 (
		.q (cell6_1Q),
		.s (cell6_1S),
		.r (cell6_1R)
);

srlt_gate cell0_2 (
		.q (cell0_2Q),
		.s (cell0_2S),
		.r (cell0_2R)
);

srlt_gate cell1_2 (
		.q (cell1_2Q),
		.s (cell1_2S),
		.r (cell1_2R)
);

srlt_gate cell2_2 (
		.q (cell2_2Q),
		.s (cell2_2S),
		.r (cell2_2R)
);

srlt_gate cell3_2 (
		.q (cell3_2Q),
		.s (cell3_2S),
		.r (cell3_2R)
);

srlt_gate cell4_2 (
		.q (cell4_2Q),
		.s (cell4_2S),
		.r (cell4_2R)
);

srlt_gate cell5_2 (
		.q (cell5_2Q),
		.s (cell5_2S),
		.r (cell5_2R)
);

srlt_gate cell6_2 (
		.q (cell6_2Q),
		.s (cell6_2S),
		.r (cell6_2R)
);

srlt_gate cell0_3 (
		.q (cell0_3Q),
		.s (cell0_3S),
		.r (cell0_3R)
);

srlt_gate cell1_3 (
		.q (cell1_3Q),
		.s (cell1_3S),
		.r (cell1_3R)
);

srlt_gate cell2_3 (
		.q (cell2_3Q),
		.s (cell2_3S),
		.r (cell2_3R)
);

srlt_gate cell3_3 (
		.q (cell3_3Q),
		.s (cell3_3S),
		.r (cell3_3R)
);

srlt_gate cell4_3 (
		.q (cell4_3Q),
		.s (cell4_3S),
		.r (cell4_3R)
);

srlt_gate cell5_3 (
		.q (cell5_3Q),
		.s (cell5_3S),
		.r (cell5_3R)
);

srlt_gate cell6_3 (
		.q (cell6_3Q),
		.s (cell6_3S),
		.r (cell6_3R)
);

srlt_gate cell0_4 (
		.q (cell0_4Q),
		.s (cell0_4S),
		.r (cell0_4R)
);

srlt_gate cell1_4 (
		.q (cell1_4Q),
		.s (cell1_4S),
		.r (cell1_4R)
);

srlt_gate cell2_4 (
		.q (cell2_4Q),
		.s (cell2_4S),
		.r (cell2_4R)
);

srlt_gate cell3_4 (
		.q (cell3_4Q),
		.s (cell3_4S),
		.r (cell3_4R)
);

srlt_gate cell4_4 (
		.q (cell4_4Q),
		.s (cell4_4S),
		.r (cell4_4R)
);

srlt_gate cell5_4 (
		.q (cell5_4Q),
		.s (cell5_4S),
		.r (cell5_4R)
);

srlt_gate cell6_4 (
		.q (cell6_4Q),
		.s (cell6_4S),
		.r (cell6_4R)
);

endmodule
